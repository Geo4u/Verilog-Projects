`timescale 1ns / 1ps
module updown_testbench();   //testbench declaration here 
reg clk, reset,up_down,pause; //inputs
reg [3:0] bin_in;
wire [6:0] hex_out;
up_down dut ( .clk(clk), .reset(reset), .up_down(up_down), .hex_out(hex_out), .pause(pause)
);
initial
begin
reset = 1'b1;#100; reset = 1'b0;#100; end
 always
6/12
begin up_down=1'b1;#400; up_down=1'b0;#1000; end
always
begin
clk = 1'b0;#10; clk = 1'b1;#10; end endmodule
 
